library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

package State_Condition is
    
    type state_type is (IDLE, SELECTMODE, GUESTIN, INPUT_USER, OVERLOAD); --masih ada pengurangan

end package;